-- Copyright (C) 2023  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 22.1std.1 Build 917 02/14/2023 SC Lite Edition"
-- CREATED		"Thu Mar 28 11:06:01 2024"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY mini_cpu IS 
	PORT
	(
		IOINBUS :  IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		KEY :  IN  STD_LOGIC_VECTOR(0 TO 0);
		SW :  IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		IOW :  OUT  STD_LOGIC;
		IOR :  OUT  STD_LOGIC;
		HEX0 :  OUT  STD_LOGIC_VECTOR(0 TO 6);
		HEX10 :  OUT  STD_LOGIC;
		HEX11 :  OUT  STD_LOGIC;
		HEX12 :  OUT  STD_LOGIC;
		HEX13 :  OUT  STD_LOGIC;
		HEX14 :  OUT  STD_LOGIC;
		HEX15 :  OUT  STD_LOGIC;
		HEX16 :  OUT  STD_LOGIC;
		HEX2 :  OUT  STD_LOGIC_VECTOR(0 TO 6);
		HEX30 :  OUT  STD_LOGIC;
		HEX31 :  OUT  STD_LOGIC;
		HEX32 :  OUT  STD_LOGIC;
		HEX33 :  OUT  STD_LOGIC;
		HEX34 :  OUT  STD_LOGIC;
		HEX35 :  OUT  STD_LOGIC;
		HEX36 :  OUT  STD_LOGIC;
		HEX4 :  OUT  STD_LOGIC_VECTOR(0 TO 6);
		HEX50 :  OUT  STD_LOGIC;
		HEX51 :  OUT  STD_LOGIC;
		HEX52 :  OUT  STD_LOGIC;
		HEX53 :  OUT  STD_LOGIC;
		HEX54 :  OUT  STD_LOGIC;
		HEX55 :  OUT  STD_LOGIC;
		HEX56 :  OUT  STD_LOGIC;
		IOADDRESS :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END mini_cpu;

ARCHITECTURE bdf_type OF mini_cpu IS 

COMPONENT reg
GENERIC (size : INTEGER
			);
	PORT(en : IN STD_LOGIC;
		 data_in : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 data_out : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT bus_mux2
GENERIC (busSize : INTEGER
			);
	PORT(sel : IN STD_LOGIC;
		 busA : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 busB : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 Q : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT bus_mux2_8b
	PORT(sel : IN STD_LOGIC;
		 busA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 busB : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 Q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT decoder
	PORT(addr : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 Q : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT bcd_to_hex
	PORT(bcd_in : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 hex_out : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END COMPONENT;

COMPONENT io_pipeline
	PORT(clk : IN STD_LOGIC;
		 en : IN STD_LOGIC;
		 reset : IN STD_LOGIC;
		 iData : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 iRegA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 op : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 opHigh : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 opLow : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 fetchE : OUT STD_LOGIC;
		 io_write : OUT STD_LOGIC;
		 io_read : OUT STD_LOGIC;
		 regA_updt : OUT STD_LOGIC;
		 oAddress : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 oData : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 oRegA : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT math_pipeline
	PORT(clk : IN STD_LOGIC;
		 en : IN STD_LOGIC;
		 reset : IN STD_LOGIC;
		 flags : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 op : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 regA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 regB : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 writeR : OUT STD_LOGIC;
		 fetchE : OUT STD_LOGIC;
		 flgUpd : OUT STD_LOGIC;
		 outFlg : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 regC : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT decoder3
	PORT(addr : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 Q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT memory_pipeline
	PORT(clk : IN STD_LOGIC;
		 en : IN STD_LOGIC;
		 reset : IN STD_LOGIC;
		 i_mem : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 i_regA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 i_regB : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 i_regC : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 op : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 opDataH : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 opDataL : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 fetchE : OUT STD_LOGIC;
		 fetchMem : OUT STD_LOGIC;
		 outAddr : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 output : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 outputPC : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 updtBus : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
	);
END COMPONENT;

COMPONENT fetcher
	PORT(clk : IN STD_LOGIC;
		 fetch_en : IN STD_LOGIC;
		 reset : IN STD_LOGIC;
		 data_in : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 pline_en : OUT STD_LOGIC;
		 pc_en : OUT STD_LOGIC;
		 op : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 operand_a : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 operand_b : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 pline_sel : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT increment_reg
GENERIC (reg_size : INTEGER
			);
	PORT(clock : IN STD_LOGIC;
		 incr_en : IN STD_LOGIC;
		 update : IN STD_LOGIC;
		 reset : IN STD_LOGIC;
		 inData : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 outData : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ram
	PORT(wren : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 address : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 data : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT rom
	PORT(clock : IN STD_LOGIC;
		 address : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	addrBus :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	AUpdate :  STD_LOGIC;
SIGNAL	DATA_OUT :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	dataA :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	dataB :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	FLAG_OUT :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	FLAG_UP :  STD_LOGIC;
SIGNAL	fm :  STD_LOGIC;
SIGNAL	HEX120 :  STD_LOGIC;
SIGNAL	HEX121 :  STD_LOGIC;
SIGNAL	HEX122 :  STD_LOGIC;
SIGNAL	HEX123 :  STD_LOGIC;
SIGNAL	HEX124 :  STD_LOGIC;
SIGNAL	HEX125 :  STD_LOGIC;
SIGNAL	HEX126 :  STD_LOGIC;
SIGNAL	HEX127 :  STD_LOGIC;
SIGNAL	HEX340 :  STD_LOGIC;
SIGNAL	HEX341 :  STD_LOGIC;
SIGNAL	HEX342 :  STD_LOGIC;
SIGNAL	HEX343 :  STD_LOGIC;
SIGNAL	HEX344 :  STD_LOGIC;
SIGNAL	HEX345 :  STD_LOGIC;
SIGNAL	HEX346 :  STD_LOGIC;
SIGNAL	HEX347 :  STD_LOGIC;
SIGNAL	HEX560 :  STD_LOGIC;
SIGNAL	HEX561 :  STD_LOGIC;
SIGNAL	HEX562 :  STD_LOGIC;
SIGNAL	HEX563 :  STD_LOGIC;
SIGNAL	HEX564 :  STD_LOGIC;
SIGNAL	HEX565 :  STD_LOGIC;
SIGNAL	HEX566 :  STD_LOGIC;
SIGNAL	HEX567 :  STD_LOGIC;
SIGNAL	io_regA :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	iow_data :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	outAddr :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	outMemPline :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	PC :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	PC_IN :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	RAM_DATA :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	regA :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	regB :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	regC :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	ROM_DATA :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	rst :  STD_LOGIC;
SIGNAL	selector :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	updtSelector :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC_VECTOR(6 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC_VECTOR(6 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC_VECTOR(6 DOWNTO 0);

SIGNAL	GDFX_TEMP_SIGNAL_8 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_7 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_6 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_5 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_4 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_3 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_2 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_1 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_0 :  STD_LOGIC_VECTOR(7 DOWNTO 0);

BEGIN 
HEX10 <= SYNTHESIZED_WIRE_47(6);
HEX11 <= SYNTHESIZED_WIRE_47(5);
HEX12 <= SYNTHESIZED_WIRE_47(4);
HEX13 <= SYNTHESIZED_WIRE_47(3);
HEX14 <= SYNTHESIZED_WIRE_47(2);
HEX15 <= SYNTHESIZED_WIRE_47(1);
HEX16 <= SYNTHESIZED_WIRE_47(0);
HEX30 <= SYNTHESIZED_WIRE_48(6);
HEX31 <= SYNTHESIZED_WIRE_48(5);
HEX32 <= SYNTHESIZED_WIRE_48(4);
HEX33 <= SYNTHESIZED_WIRE_48(3);
HEX34 <= SYNTHESIZED_WIRE_48(2);
HEX35 <= SYNTHESIZED_WIRE_48(1);
HEX36 <= SYNTHESIZED_WIRE_48(0);
HEX50 <= SYNTHESIZED_WIRE_49(6);
HEX51 <= SYNTHESIZED_WIRE_49(5);
HEX52 <= SYNTHESIZED_WIRE_49(4);
HEX53 <= SYNTHESIZED_WIRE_49(3);
HEX54 <= SYNTHESIZED_WIRE_49(2);
HEX55 <= SYNTHESIZED_WIRE_49(1);
HEX56 <= SYNTHESIZED_WIRE_49(0);

GDFX_TEMP_SIGNAL_8 <= (HEX567 & HEX566 & HEX565 & HEX564);
GDFX_TEMP_SIGNAL_7 <= (HEX563 & HEX562 & HEX561 & HEX560);
GDFX_TEMP_SIGNAL_6 <= (HEX347 & HEX346 & HEX345 & HEX344);
GDFX_TEMP_SIGNAL_5 <= (HEX343 & HEX342 & HEX341 & HEX340);
GDFX_TEMP_SIGNAL_4 <= (HEX127 & HEX126 & HEX125 & HEX124);
GDFX_TEMP_SIGNAL_3 <= (HEX123 & HEX122 & HEX121 & HEX120);
HEX567 <= GDFX_TEMP_SIGNAL_2(7);
HEX566 <= GDFX_TEMP_SIGNAL_2(6);
HEX565 <= GDFX_TEMP_SIGNAL_2(5);
HEX564 <= GDFX_TEMP_SIGNAL_2(4);
HEX563 <= GDFX_TEMP_SIGNAL_2(3);
HEX562 <= GDFX_TEMP_SIGNAL_2(2);
HEX561 <= GDFX_TEMP_SIGNAL_2(1);
HEX560 <= GDFX_TEMP_SIGNAL_2(0);

HEX347 <= GDFX_TEMP_SIGNAL_1(7);
HEX346 <= GDFX_TEMP_SIGNAL_1(6);
HEX345 <= GDFX_TEMP_SIGNAL_1(5);
HEX344 <= GDFX_TEMP_SIGNAL_1(4);
HEX343 <= GDFX_TEMP_SIGNAL_1(3);
HEX342 <= GDFX_TEMP_SIGNAL_1(2);
HEX341 <= GDFX_TEMP_SIGNAL_1(1);
HEX340 <= GDFX_TEMP_SIGNAL_1(0);

HEX127 <= GDFX_TEMP_SIGNAL_0(7);
HEX126 <= GDFX_TEMP_SIGNAL_0(6);
HEX125 <= GDFX_TEMP_SIGNAL_0(5);
HEX124 <= GDFX_TEMP_SIGNAL_0(4);
HEX123 <= GDFX_TEMP_SIGNAL_0(3);
HEX122 <= GDFX_TEMP_SIGNAL_0(2);
HEX121 <= GDFX_TEMP_SIGNAL_0(1);
HEX120 <= GDFX_TEMP_SIGNAL_0(0);



b2v_A_Register : reg
GENERIC MAP(size => 8
			)
PORT MAP(en => SYNTHESIZED_WIRE_0,
		 data_in => SYNTHESIZED_WIRE_1,
		 data_out => regA);


b2v_addrMux : bus_mux2
GENERIC MAP(busSize => 16
			)
PORT MAP(sel => fm,
		 busA => PC,
		 busB => outAddr,
		 Q => addrBus);


b2v_B_Register : reg
GENERIC MAP(size => 8
			)
PORT MAP(en => updtSelector(2),
		 data_in => SYNTHESIZED_WIRE_44,
		 data_out => regB);


b2v_C_Register : reg
GENERIC MAP(size => 8
			)
PORT MAP(en => SYNTHESIZED_WIRE_3,
		 data_in => SYNTHESIZED_WIRE_44,
		 data_out => regC);


b2v_dataMux : bus_mux2_8b
PORT MAP(sel => SYNTHESIZED_WIRE_5,
		 busA => RAM_DATA,
		 busB => ROM_DATA,
		 Q => DATA_OUT);


b2v_dbg_muxA : bus_mux2_8b
PORT MAP(sel => SW(1),
		 busA => PC(7 DOWNTO 0),
		 busB => regA,
		 Q => GDFX_TEMP_SIGNAL_0);


b2v_dbg_muxB : bus_mux2_8b
PORT MAP(sel => SW(1),
		 busA => PC(15 DOWNTO 8),
		 busB => regB,
		 Q => GDFX_TEMP_SIGNAL_1);


b2v_dbg_muxC : bus_mux2_8b
PORT MAP(sel => SW(1),
		 busA => DATA_OUT,
		 busB => regC,
		 Q => GDFX_TEMP_SIGNAL_2);


b2v_decode_pline_selector : decoder
PORT MAP(addr => SYNTHESIZED_WIRE_6,
		 Q => selector);


SYNTHESIZED_WIRE_24 <= SYNTHESIZED_WIRE_7 OR SYNTHESIZED_WIRE_8 OR SYNTHESIZED_WIRE_9;


b2v_FLAGS : reg
GENERIC MAP(size => 8
			)
PORT MAP(en => FLAG_UP,
		 data_in => FLAG_OUT,
		 data_out => SYNTHESIZED_WIRE_19);


b2v_hexA : bcd_to_hex
PORT MAP(bcd_in => GDFX_TEMP_SIGNAL_3,
		 hex_out => HEX0);


b2v_hexB : bcd_to_hex
PORT MAP(bcd_in => GDFX_TEMP_SIGNAL_4,
		 hex_out => SYNTHESIZED_WIRE_47);


b2v_hexC : bcd_to_hex
PORT MAP(bcd_in => GDFX_TEMP_SIGNAL_5,
		 hex_out => HEX2);


b2v_hexD : bcd_to_hex
PORT MAP(bcd_in => GDFX_TEMP_SIGNAL_6,
		 hex_out => SYNTHESIZED_WIRE_48);


b2v_hexE : bcd_to_hex
PORT MAP(bcd_in => GDFX_TEMP_SIGNAL_7,
		 hex_out => HEX4);


b2v_hexF : bcd_to_hex
PORT MAP(bcd_in => GDFX_TEMP_SIGNAL_8,
		 hex_out => SYNTHESIZED_WIRE_49);


SYNTHESIZED_WIRE_18 <= SYNTHESIZED_WIRE_45 AND selector(1);


SYNTHESIZED_WIRE_5 <= NOT(addrBus(15));



SYNTHESIZED_WIRE_22 <= SYNTHESIZED_WIRE_45 AND selector(2);


SYNTHESIZED_WIRE_44 <= outMemPline OR SYNTHESIZED_WIRE_12;


SYNTHESIZED_WIRE_16 <= SYNTHESIZED_WIRE_45 AND selector(3);


SYNTHESIZED_WIRE_3 <= updtSelector(3) OR SYNTHESIZED_WIRE_14;


SYNTHESIZED_WIRE_0 <= AUpdate OR updtSelector(1);


SYNTHESIZED_WIRE_1 <= io_regA OR SYNTHESIZED_WIRE_44;


b2v_io_pline : io_pipeline
PORT MAP(clk => SW(0),
		 en => SYNTHESIZED_WIRE_16,
		 reset => rst,
		 iData => IOINBUS,
		 iRegA => regA,
		 op => SYNTHESIZED_WIRE_46,
		 opHigh => dataB,
		 opLow => dataA,
		 fetchE => SYNTHESIZED_WIRE_8,
		 io_write => IOW,
		 io_read => IOR,
		 regA_updt => AUpdate,
		 oAddress => IOADDRESS,
		 oRegA => io_regA);


b2v_math_pline : math_pipeline
PORT MAP(clk => SW(0),
		 en => SYNTHESIZED_WIRE_18,
		 reset => rst,
		 flags => SYNTHESIZED_WIRE_19,
		 op => SYNTHESIZED_WIRE_46,
		 regA => regA,
		 regB => regB,
		 writeR => SYNTHESIZED_WIRE_14,
		 fetchE => SYNTHESIZED_WIRE_9,
		 flgUpd => FLAG_UP,
		 outFlg => FLAG_OUT,
		 regC => SYNTHESIZED_WIRE_12);


b2v_memdecode : decoder3
PORT MAP(addr => SYNTHESIZED_WIRE_21,
		 Q => updtSelector);


b2v_memory_pline : memory_pipeline
PORT MAP(clk => SW(0),
		 en => SYNTHESIZED_WIRE_22,
		 reset => rst,
		 i_mem => DATA_OUT,
		 i_regA => regA,
		 i_regB => regB,
		 i_regC => regC,
		 op => SYNTHESIZED_WIRE_46,
		 opDataH => dataB,
		 opDataL => dataA,
		 fetchE => SYNTHESIZED_WIRE_7,
		 fetchMem => fm,
		 outAddr => outAddr,
		 output => outMemPline,
		 outputPC => PC_IN,
		 updtBus => SYNTHESIZED_WIRE_21);


b2v_op_fetcher : fetcher
PORT MAP(clk => SW(0),
		 fetch_en => SYNTHESIZED_WIRE_24,
		 reset => rst,
		 data_in => DATA_OUT,
		 pline_en => SYNTHESIZED_WIRE_45,
		 pc_en => SYNTHESIZED_WIRE_25,
		 op => SYNTHESIZED_WIRE_46,
		 operand_a => dataA,
		 operand_b => dataB,
		 pline_sel => SYNTHESIZED_WIRE_6);


b2v_program_counter : increment_reg
GENERIC MAP(reg_size => 16
			)
PORT MAP(clock => SW(0),
		 incr_en => SYNTHESIZED_WIRE_25,
		 update => updtSelector(4),
		 reset => rst,
		 inData => PC_IN,
		 outData => PC);


b2v_ram_block : ram
PORT MAP(wren => updtSelector(5),
		 clock => SW(0),
		 address => addrBus,
		 data => outMemPline,
		 q => RAM_DATA);


b2v_rom_block : rom
PORT MAP(clock => SW(0),
		 address => addrBus,
		 q => ROM_DATA);

rst <= KEY(0);

HEX120 <= GDFX_TEMP_SIGNAL_0(0);
HEX121 <= GDFX_TEMP_SIGNAL_0(1);
HEX122 <= GDFX_TEMP_SIGNAL_0(2);
HEX123 <= GDFX_TEMP_SIGNAL_0(3);
HEX124 <= GDFX_TEMP_SIGNAL_0(4);
HEX125 <= GDFX_TEMP_SIGNAL_0(5);
HEX126 <= GDFX_TEMP_SIGNAL_0(6);
HEX127 <= GDFX_TEMP_SIGNAL_0(7);
HEX340 <= GDFX_TEMP_SIGNAL_1(0);
HEX341 <= GDFX_TEMP_SIGNAL_1(1);
HEX342 <= GDFX_TEMP_SIGNAL_1(2);
HEX343 <= GDFX_TEMP_SIGNAL_1(3);
HEX344 <= GDFX_TEMP_SIGNAL_1(4);
HEX345 <= GDFX_TEMP_SIGNAL_1(5);
HEX346 <= GDFX_TEMP_SIGNAL_1(6);
HEX347 <= GDFX_TEMP_SIGNAL_1(7);
HEX560 <= GDFX_TEMP_SIGNAL_2(0);
HEX561 <= GDFX_TEMP_SIGNAL_2(1);
HEX562 <= GDFX_TEMP_SIGNAL_2(2);
HEX563 <= GDFX_TEMP_SIGNAL_2(3);
HEX564 <= GDFX_TEMP_SIGNAL_2(4);
HEX565 <= GDFX_TEMP_SIGNAL_2(5);
HEX566 <= GDFX_TEMP_SIGNAL_2(6);
HEX567 <= GDFX_TEMP_SIGNAL_2(7);
END bdf_type;